module tf_ROM 
    #(parameter addr_rom_width = 6,
                 data_width = 36,
                 depth_rom = 40)
    (
    input clk,
    input [addr_rom_width-1:0] A,
    input IREN,
    output reg [data_width-1:0] Q);
    
    always@(posedge clk)
    begin
    if(IREN == 1'b1) begin
    case(A)
    9'd0:  Q <= 36'b011011111001111010100011101000111111;
    9'd1:  Q <= 36'b001101110101101010101110100010100110;
    9'd2:  Q <= 36'b101001100100110101100110100010001001;
    9'd3:  Q <= 36'b100110000100000000101101001001011011;
    9'd4:  Q <= 36'b001100011110110111111101101100100111;
    9'd5:  Q <= 36'b001001000011110111010010110000110000;
    9'd6:  Q <= 36'b100011100000001001011100000010010000;
    9'd7:  Q <= 36'b101100010001100010100100111110110000;
    9'd8:  Q <= 36'b010011110111101011000100110000101110;
    9'd9:  Q <= 36'b001100000100110101100110000010001110;
    9'd10: Q <= 36'b100100011011100100111001111110101101;
    9'd11: Q <= 36'b011111001000010111100001001010101011;
    9'd12: Q <= 36'b100100000101100101101100010000001110;
    9'd13: Q <= 36'b010010111011101011011100111010111101;
    9'd14: Q <= 36'b010010110001011001000100001101111101;
    9'd15: Q <= 36'b100011110000101001000110001010110100;
    9'd16: Q <= 36'b101011110110111001010100100100011001;
    9'd17: Q <= 36'b101011011010001000110000000110001111;
    9'd18: Q <= 36'b101111011101010111001000111110001000;
    9'd19: Q <= 36'b101001100111100110010111000001110100;
    9'd20: Q <= 36'b011101111111100001010100011100010000;
    9'd21: Q <= 36'b001001011000010001001110110000100001;
    9'd22: Q <= 36'b000001100001100100100001100010111111;
    9'd23: Q <= 36'b011100000101000100010010010001110011;
    9'd24: Q <= 36'b100001000010000110011000011000000010;
    9'd25: Q <= 36'b000011111110010001111101110101110001;
    9'd26: Q <= 36'b000000000110110000101101100101110011;
    9'd27: Q <= 36'b000110011000001000110010100000101001;
    9'd28: Q <= 36'b100001010011100011001010100101101110;
    9'd29: Q <= 36'b000001011000100010010111101010101001;
    9'd30: Q <= 36'b010011100101000001011001010001001101;
    9'd31: Q <= 36'b100100101000010000010100111010100100;
    9'd32: Q <= 36'b001011001010110001101010000001101101;
    9'd33: Q <= 36'b000110000000010010110100000100111111;
    9'd34: Q <= 36'b100101100010110111000001110101111011;
    9'd35: Q <= 36'b010010011010100011001101010010001011;
    9'd36: Q <= 36'b010011100110111001111101100010011110;
    9'd37: Q <= 36'b001000011101101001001110011100001111;
    9'd38: Q <= 36'b101111011000010000111111111010000101;
    9'd39: Q <= 36'b101111100100000000011110000001110000;
    9'd40: Q <= 42'b101111111111100000000000100110111111;
    9'd41: Q <= 42'b001101001001001010010111100000000110;
    9'd42: Q <= 42'b100100111000100110110010111000000110;
    endcase end         
    end
endmodule